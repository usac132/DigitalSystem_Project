module print_score_7seg(

)
// score을 7segment display에 표시

// 기존에 만들었던거 그냥 갖다 쓰면 될듯

endmodule