module print_score_7seg(
    input [6:0] score,
    output //7segment control, display
);
// score을 7segment display에 표시

// 기존에 수업때 만들었던거 수정해서 갖다 넣기

endmodule